// frame_controller.v
// CMPE 670 Project Fall 2023
// Author(s):
//  John Evans
module frame_controller (
    // clock and control
    input        i_clk,
    input        i_rst,
    input        i_row_cnt,
    input        i_col_cnt,
    //
    input        i_pyld_data_valid,
    input        i_line_fifo_ready,
    // outputs
    output       o_data_req
);





endmodule