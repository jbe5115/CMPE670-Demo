// fpc.v
// CMPE 670 Project Fall 2023
// Author(s):
//   
module fpc (
    // clock and control
    input        i_clk,
    input        i_rst,

    input        i_pyld_data_valid,

    output       o_row_cnt,
    output       o_col_cnt
);


endmodule